// Created by prof. Mingu Kang @VVIP Lab in UCSD ECE department
// Please do not spread this code without permission 
module ofifo (clk, in, out, rd, wr, o_full, reset, o_ready, o_valid);

  parameter col  = 8;
  parameter psum_bw = 16;

  input  clk;
  input  [col - 1 : 0] wr;
  input  rd;
  input  reset;
  input  [psum_bw * col - 1 : 0] in;
  output [psum_bw * col - 1 : 0] out;
  output o_full;
  output o_ready;
  output o_valid;

  wire [col - 1 : 0] empty;
  wire [col - 1 : 0] full;
  reg  rd_en;
  
  genvar i;

  assign o_ready = !(|full);
  assign o_full  = (|full);
  assign o_valid = !(|empty);

  generate
	  for (i=0; i<col ; i=i+1) begin : col_num
			fifo_depth36 #(.bw(psum_bw)) fifo_instance (
			  .rd_clk(clk),
			  .wr_clk(clk),
			  .rd(rd_en),
			  .wr(wr[i]),
			  .reset(reset),
			  .o_full(full[i]),
			  .o_empty(empty[i]),
			  .in(in[(i+1)*psum_bw - 1 : i*psum_bw]),
			  .out(out[(i+1)*psum_bw - 1 : i*psum_bw])
			  );
	  end
	endgenerate

  always @ (posedge clk) begin
   if (reset) begin
      rd_en <= 0;
   end
   else begin
      rd_en <= rd;
   end
 
  end


 

endmodule
